library verilog;
use verilog.vl_types.all;
entity macrofunction_vlg_vec_tst is
end macrofunction_vlg_vec_tst;
