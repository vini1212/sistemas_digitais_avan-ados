library verilog;
use verilog.vl_types.all;
entity Lookahead_vlg_vec_tst is
end Lookahead_vlg_vec_tst;
