library verilog;
use verilog.vl_types.all;
entity RippleCarry_vlg_vec_tst is
end RippleCarry_vlg_vec_tst;
